-- Memory controller generated from the DSP toolbox
-- Electronics Systems, http://www.es.isy.liu.se/

library ieee;
use ieee.std_logic_1164.all;

entity memorycontroller2 is
port(
state : in integer range 0 to 47;
adress : out integer range 0 to 9;
enable, readwrite : out std_logic);
end memorycontroller2;

architecture generated of memorycontroller2 is
begin
with state select
adress <= 
1 when 0,
0 when 1,
5 when 2,
1 when 3,
2 when 4,
2 when 5,
9 when 6,
3 when 7,
6 when 8,
4 when 9,
4 when 10,
4 when 11,
8 when 12,
5 when 13,
2 when 14,
2 when 15,
5 when 16,
5 when 17,
0 when 18,
0 when 19,
0 when 20,
0 when 21,
0 when 22,
6 when 23,
2 when 24,
0 when 25,
7 when 26,
2 when 27,
7 when 29,
8 when 31,
2 when 32,
2 when 33,
2 when 34,
2 when 35,
1 when 36,
9 when 37,
7 when 38,
1 when 39,
3 when 40,
7 when 41,
0 when 42,
4 when 44,
8 when 46,
8 when 47,
0 when others;

with state select
readwrite <= 
'1' when 0,
'0' when 1,
'1' when 2,
'0' when 3,
'1' when 4,
'0' when 5,
'1' when 6,
'0' when 7,
'1' when 8,
'0' when 9,
'1' when 10,
'0' when 11,
'1' when 12,
'0' when 13,
'1' when 14,
'0' when 15,
'1' when 16,
'0' when 17,
'1' when 18,
'0' when 19,
'1' when 20,
'0' when 21,
'1' when 22,
'0' when 23,
'1' when 24,
'0' when 25,
'1' when 26,
'0' when 27,
'0' when 29,
'0' when 31,
'1' when 32,
'0' when 33,
'1' when 34,
'0' when 35,
'1' when 36,
'0' when 37,
'1' when 38,
'0' when 39,
'1' when 40,
'0' when 41,
'1' when 42,
'1' when 44,
'1' when 46,
'0' when 47,
'-' when others;

with state select
enable <= 
'1' when 0,
'1' when 1,
'1' when 2,
'1' when 3,
'1' when 4,
'1' when 5,
'1' when 6,
'1' when 7,
'1' when 8,
'1' when 9,
'1' when 10,
'1' when 11,
'1' when 12,
'1' when 13,
'1' when 14,
'1' when 15,
'1' when 16,
'1' when 17,
'1' when 18,
'1' when 19,
'1' when 20,
'1' when 21,
'1' when 22,
'1' when 23,
'1' when 24,
'1' when 25,
'1' when 26,
'1' when 27,
'1' when 29,
'1' when 31,
'1' when 32,
'1' when 33,
'1' when 34,
'1' when 35,
'1' when 36,
'1' when 37,
'1' when 38,
'1' when 39,
'1' when 40,
'1' when 41,
'1' when 42,
'1' when 44,
'1' when 46,
'1' when 47,
'0' when others;

end generated;
